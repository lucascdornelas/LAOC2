library verilog;
use verilog.vl_types.all;
entity parte1maq2 is
    port(
        clock           : in     vl_logic;
        SW              : in     vl_logic_vector(1 downto 0)
    );
end parte1maq2;
