
module pratica_3_tomasulo(
	input clock
);
	CDB cdb (clock);
endmodule