library verilog;
use verilog.vl_types.all;
entity pratica_3_tomasulo is
    port(
        clock           : in     vl_logic;
        Reset           : in     vl_logic;
        Run             : in     vl_logic
    );
end pratica_3_tomasulo;
